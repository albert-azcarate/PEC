LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY L1_T3 IS
	 PORT( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
	 LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END L1_T3;
ARCHITECTURE Structure OF L1_T3 IS
BEGIN
			LEDR<=SW;
END Structure; 
