-- 
-- Input: ->  bits
-- Output: ->  bits

LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY NOM IS

-- generics


-- ports
	PORT(	
			);
			
END NOM;

ARCHITECTURE Structure OF NOM IS

-- constants

-- components

-- variables

BEGIN
	
	-- mapping
	
	
END Structure;